`timescale 1ns / 1ps
module spi(
	input rst, clk, newd,
  input [11:0]din,
  output reg mosi,
  output reg cs, sclk
);
  
  int countc = 0;
  int count = 0;
  
  typedef enum bit[1:0]{idle = 2'b00, send = 2'b01}state_type;
  state_type state = idle;
  
  
  ///sclk generation
  always@(posedge clk)begin
    if(rst == 1'b1) begin countc <= 0; sclk <= 1'b0;end
    else begin
      if(countc < 10) countc <= countc + 1;
      else begin
        countc <= 0;
        sclk <= ~sclk;
      end
    end
  end
  

  reg [11:0]temp;
  
  always@(posedge sclk)begin
    
    if(rst == 1'b1)begin
      cs <= 1'b1;
      mosi <= 1'b0;
    end
    
    else begin
      case(state)
        
        idle:begin
          if(newd == 1'b1)begin
            cs <= 1'b0;
            temp <= din;
            state <= send;
          end
          else begin
            state <= idle;
            temp <= 8'h00;
          end
        end
        
        send:begin
          
          if(count < 12)begin
            mosi <= temp[count];
            count <= count + 1;
           end
          else begin
            count <= 0;
            cs <= 1'b1;
            mosi <= 1'b0;
            state <= idle;
          end
          
        end
        
        default: state<=idle;
        
      endcase
    end///-
    
  end//-
  
endmodule
interface spi_if;
  logic rst, clk, newd;
  logic [11:0]din;
  logic mosi,cs, sclk;
endinterface